  
 --******************************************************************************************
 --*  COMPANY    :  Microsoft                                                               *
 --*  NAME       :  ece                                                                     *
 --*  BOARD      :  ProceV_D8                                                               *
 --*  IC#        :  1                                                                       *
 --*  Created    :  Sat Aug 12 20:18:15 2017                                                *
 --*  This file  was  generated by  ProcWizard Application  version 9.5.0.0                 *
 --*  Copyright (C) 2017. All Rights Reserved to Gidel Ltd                                  *
 --******************************************************************************************
  
  
  
  
  
 LIBRARY   ieee;
 USE       ieee.std_logic_1164.all;
 USE       ieee.std_logic_unsigned.all;
 


 PACKAGE dma_package IS
   TYPE   arr_19x0_31x0     IS ARRAY  ( 19 DOWNTO 0 )  OF   STD_LOGIC_VECTOR( 31 DOWNTO 0 );
   TYPE   arr_2x0_31x0      IS ARRAY  ( 2  DOWNTO 0 )  OF   STD_LOGIC_VECTOR( 31 DOWNTO 0 );
   TYPE   arr_39x0_31x0     IS ARRAY  ( 39 DOWNTO 0 )  OF   STD_LOGIC_VECTOR( 31 DOWNTO 0 );
 END dma_package;
  
 --======================================================================
 --=                   Use Altera Libraries For VHDL                    =
 --======================================================================
 LIBRARY altera;
 USE altera.altera_primitives_components.all;
  
  
 LIBRARY   ieee;
 USE       ieee.std_logic_1164.all;
 USE       ieee.std_logic_unsigned.all;
 USE       ieee.std_logic_arith.all;
   
   
 LIBRARY   work;
 USE       work.dma_package.all;
  
 ENTITY   dma   IS
     PORT(
 --======================================================================
 --=                         Clocks & Globals                           =
 --======================================================================
  ref_clk                        : IN    STD_LOGIC;                          -- 25 MHz reference clock input pin
  mem_ref_clk                    : IN    STD_LOGIC;                          -- 125MHz, memory reference clock input pin
  ext_clk                        : IN    STD_LOGIC;                          -- User external clock from SMA
  ext_resetn                     : IN    STD_LOGIC;                          -- Used in stand-alone from push button
  scl                            : INOUT STD_LOGIC;                          -- SODIMM Serial clock. Used to synchronize communication to and from the I2C bus
  sda                            : INOUT STD_LOGIC;                          -- SODIMM Serial data:  Used to transfer addresses and data into and out of the I2C bus
  ledn                           : OUT   STD_LOGIC_VECTOR( 4  DOWNTO 1 );    -- General Purpose User LEDs; 0: light on
  status_ledn                    : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 1 );    -- Status LEDs; 0: light on
  g_reserved                     : INOUT STD_LOGIC_VECTOR( 33 DOWNTO 0 );    -- Gidel reserved IO bus
  
 --======================================================================
 --=                       PCIe Bus Connections                         =
 --======================================================================
  pcie_refclk                    : IN    STD_LOGIC;                          -- Reference clock for the Stratix V Hard IP for PCI Express
  pcie_perst                     : IN    STD_LOGIC;                          -- Active low reset from the PCIe reset pin of the device
  pcie_rx                        : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Receive inputs. These signals are the serial inputs of lanes 7�0
  pcie_tx                        : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Transmit outputs. These signals are the serial outputs of lanes 7�0
  
 --======================================================================
 --=                    DDR3 SDRAM block B (SODIMM)                     =
 --======================================================================
  addr_b                         : OUT   STD_LOGIC_VECTOR( 15 DOWNTO 0 );    -- Address bus
  ba_b                           : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- Bank address select
  cas_b                          : OUT   STD_LOGIC;                          -- Command output(CAS) - active LOW
  cke_b                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock enable - active HIGH
  ck_b                           : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock: Differential clock outputs (positive)
  ckn_b                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock: Differential clock outputs (negative)
  cs_b                           : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Chip select - active LOW
  dq_b                           : INOUT STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Data bus
  dqm_b                          : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data mask,is an output mask signal for write data (byte enable)
  dqs_b                          : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data strobe: Differential data strobes (positive)
  dqsn_b                         : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data strobe: Differential data strobes (negative)
  we_b                           : OUT   STD_LOGIC;                          -- Write enable - active LOW
  ras_b                          : OUT   STD_LOGIC;                          -- Command output(RAS) - active LOW
  odt_b                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- On-die termination enable - active HIGH
  resetn_b                       : OUT   STD_LOGIC;                          -- asynchronous SODIMM Reset - active LOW
  event_b                        : IN    STD_LOGIC;                          -- 1: SODIMM critical temperature thresholds have been exceeded
  rzq_b                          : IN    STD_LOGIC;                          -- Used for OCT calibration, the RZQ pin is connected to GND through an external 240-Ohm reference resistor
  
 --======================================================================
 --=                    DDR3 SDRAM block C (SODIMM)                     =
 --======================================================================
  addr_c                         : OUT   STD_LOGIC_VECTOR( 15 DOWNTO 0 );    -- Address bus
  ba_c                           : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- Bank address select
  cas_c                          : OUT   STD_LOGIC;                          -- Command output(CAS) - active LOW
  cke_c                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock enable - active HIGH
  ck_c                           : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock: Differential clock outputs (positive)
  ckn_c                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock: Differential clock outputs (negative)
  cs_c                           : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Chip select - active LOW
  dq_c                           : INOUT STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Data bus
  dqm_c                          : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data mask,is an output mask signal for write data (byte enable)
  dqs_c                          : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data strobe: Differential data strobes (positive)
  dqsn_c                         : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Data strobe: Differential data strobes (negative)
  we_c                           : OUT   STD_LOGIC;                          -- Write enable - active LOW
  ras_c                          : OUT   STD_LOGIC;                          -- Command output(RAS) - active LOW
  odt_c                          : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- On-die termination enable - active HIGH
  resetn_c                       : OUT   STD_LOGIC;                          -- asynchronous SODIMM Reset - active LOW
  event_c                        : IN    STD_LOGIC;                          -- 1: SODIMM critical temperature thresholds have been exceeded
  rzq_c                          : IN    STD_LOGIC;                          -- Used for OCT calibration, the RZQ pin is connected to GND through an external 240-Ohm reference resistor
  
 --======================================================================
 --=                    DDR2 SRAM block D (Onboard)                     =
 --======================================================================
  dq_d                           : INOUT STD_LOGIC_VECTOR( 35 DOWNTO 0 );    -- Data bus
  ldn_d                          : OUT   STD_LOGIC;                          -- Synchronous load - active LOW
  bwsn_d                         : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 0 );    -- Byte Write Select - active LOW
  r_wn_d                         : OUT   STD_LOGIC;                          -- 1: Synchronous read 0: Synchronous write
  k_d                            : OUT   STD_LOGIC;                          -- Positive output clock input
  cq_d                           : IN    STD_LOGIC;                          -- Clock (positive) synchronized to the input data
  cqn_d                          : IN    STD_LOGIC;                          -- Do not use
  qvld_d                         : IN    STD_LOGIC;                          -- 1: valid input data. QVLD is edge aligned with CQ and CQn.
  addr_d                         : OUT   STD_LOGIC_VECTOR( 21 DOWNTO 0 );    -- Address bus
  
 --======================================================================
 --=                    DDR2 SRAM block E (Onboard)                     =
 --======================================================================
  dq_e                           : INOUT STD_LOGIC_VECTOR( 35 DOWNTO 0 );    -- Data bus
  ldn_e                          : OUT   STD_LOGIC;                          -- Synchronous load - active LOW
  bwsn_e                         : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 0 );    -- Byte Write Select - active LOW
  r_wn_e                         : OUT   STD_LOGIC;                          -- 1: Synchronous read 0: Synchronous write
  k_e                            : OUT   STD_LOGIC;                          -- Positive output clock input
  cq_e                           : IN    STD_LOGIC;                          -- Clock (positive) synchronized to the input data
  cqn_e                          : IN    STD_LOGIC;                          -- Do not use
  qvld_e                         : IN    STD_LOGIC;                          -- 1: valid input data. QVLD is edge aligned with CQ and CQn.
  addr_e                         : OUT   STD_LOGIC_VECTOR( 21 DOWNTO 0 );    -- Address bus
  
 --======================================================================
 --=                       User Buses / Signals                         =
 --======================================================================
 --======================================================================
 --=            1G PHY I/O's (Connections to on board PHY)              =
 --======================================================================
  phy_mdio                       : INOUT STD_LOGIC;                          -- Is a management data
  phy_mdc                        : OUT   STD_LOGIC;                          -- Is a management data clock reference
  phy_resetn                     : OUT   STD_LOGIC;                          -- Is a hardware reset - active LOW
  phy_rx_ctrl                    : IN    STD_LOGIC;                          -- Is a RGMII receive control
  phy_rx_clk                     : IN    STD_LOGIC;                          -- Is a RGMII receive clock
  phy_rxd                        : IN    STD_LOGIC_VECTOR( 3  DOWNTO 0 );    -- Is a RGMII receive data
  phy_tx_ctrl                    : OUT   STD_LOGIC;                          -- Is a RGMII transmit control
  phy_tx_clk                     : OUT   STD_LOGIC;                          -- Is a RGMII transmit clock
  phy_txd                        : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 0 );    -- Is a RGMII transmit data
  
 --======================================================================
 --=                               SFP A                                =
 --======================================================================
  sfp_mod_abs_a                  : IN    STD_LOGIC;                          -- 0: Module Absent, 1: Module inserted
  sfp_link_ledn_a                : OUT   STD_LOGIC;                          -- 0: led on
  sfp_trafic_ledn_a              : OUT   STD_LOGIC;                          -- 0: led on
 --======================================================================
 --=                               SFP B                                =
 --======================================================================
  sfp_mod_abs_b                  : IN    STD_LOGIC;                          -- 0: Module Absent, 1: Module inserted
  sfp_link_ledn_b                : OUT   STD_LOGIC;                          -- 0: led on
  sfp_trafic_ledn_b              : OUT   STD_LOGIC;                          -- 0: led on
  
 --======================================================================
 --=                                CXP                                 =
 --======================================================================
  cxp_prsnt_l                    : IN    STD_LOGIC;                          -- Is used to indicate when the module is plugged into the host receptacle
 --======================================================================
 --=       High Speed (HS-B) - 8 lanes transceivers connections         =
 --======================================================================
  hs_prsnt_b                     : IN    STD_LOGIC;                          -- 0: This port is connected
 --======================================================================
 --=       High Speed (HS-C) - 4 lanes transceivers connections         =
 --======================================================================
  hs_prsnt_c                     : IN    STD_LOGIC;                          -- 0: This port is connected
 --======================================================================
 --=                   External(J3) connector I/O's                     =
 --======================================================================
  j3_ext_io                      : INOUT STD_LOGIC_VECTOR( 11 DOWNTO 0 );    -- General-purpose I/O bus
  j3_ext_io_dir                  : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Bit-0 sets direction for ext_io[7:0] and bit-1 for ext_io[11:8]. (ext_io_dir=0: Inputs, ext_io_dir=1: Outputs)
 --======================================================================
 --=                       L(J4) connector I/O's                        =
 --======================================================================
  l                              : INOUT STD_LOGIC_VECTOR( 84 DOWNTO 0 );    -- Bidirectional Left bus
  l_in                           : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Left input bus
  l_io                           : INOUT STD_LOGIC_VECTOR( 19 DOWNTO 0 );    -- Left io bus
  clk_out                        : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 )     -- Clock output
     );
 END   dma;
  
  
 ARCHITECTURE  dma_arch  OF  dma  IS
 CONSTANT    RBF_VERSION_VAL                       :STD_LOGIC_VECTOR := "00000001";
  
 COMPONENT   dma_if
     PORT(
  
 --Clocks & Globals
  ref_clk                        : IN    STD_LOGIC;                          -- 25 MHz reference clock input pin
  clk0                           : OUT   STD_LOGIC;                          -- Main system clock, the max frequency is 300 MHZ
  clk                            : OUT   STD_LOGIC;                          -- User clock, the frequency is twice/triply the frequency of clk0
  clk2                           : OUT   STD_LOGIC;                          -- Is an auxiliary clock that may be used as a slow emulation clock
  mem_ref_clk_int                : OUT   STD_LOGIC;                          -- Is an internal (from PLL) memory reference clock (125MHz)
  scl                            : INOUT STD_LOGIC;                          -- Serial clock. Used to synchronize communication to and from the I2C bus
  sda                            : INOUT STD_LOGIC;                          -- Serial data: Used to transfer addresses and data into and out of the I2C bus
  status_ledn                    : OUT   STD_LOGIC_VECTOR( 3  DOWNTO 1 );    -- Status LEDs; 0: light on
  id                             : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- FPGA number identification
  g_reserved                     : INOUT STD_LOGIC_VECTOR( 33 DOWNTO 0 );    -- Gidel reserved IO bus
  g_reserved_control             : OUT   STD_LOGIC_VECTOR( 99 DOWNTO 0 );    -- Gidel reserved control bus (out)
  
 --PCIe connection
  pcie_refclk                    : IN    STD_LOGIC;                          -- Reference clock for the Hard IP for PCI Express
  pcie_perst                     : IN    STD_LOGIC;                          -- Active low reset from the PCIe reset pin of the device
  pcie_rx                        : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Receive inputs. These signals are the serial inputs of lanes 7�0
  pcie_tx                        : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- Transmit outputs. These signals are the serial outputs of lanes 7�0
  
 --Internal Bus Interface Signals
  clrn                           : OUT   STD_LOGIC;                          -- User Global Clear   (0: clear all)
  lclk                           : OUT   STD_LOGIC;                          -- Local Bus Clock
  l_wr                           : OUT   STD_LOGIC;                          -- User Write Signal (1:write)
  addr_wr                        : OUT   STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- local bus address for write operations (including burst auto address increment)
  l_data_wr                      : OUT   STD_LOGIC_VECTOR( 255 DOWNTO 0 );   -- user input local data bus
  mem_ready_wr                   : IN    STD_LOGIC;                          -- 1: end of data write transfer (memory data is valid) on rising edge of lclk
  l_rd                           : OUT   STD_LOGIC;                          -- User Read Signal (0:read)
  addr_rd                        : OUT   STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- local bus address for read operations (including burst auto address increment)
  l_data_rd                      : IN    STD_LOGIC_VECTOR( 255 DOWNTO 0 );   -- data to read back from device memories
  mem_ready_rd                   : IN    STD_LOGIC;                          -- 1: end of data read transfer (memory data is valid) on rising edge of lclk
  
 --Interrupt Logic
  interrupt                      : IN    STD_LOGIC;                          -- User interrupt
  interrupt_ack                  : OUT   STD_LOGIC;                          -- User interrupt acknowledge
  
 --DREQ Logic
  user_dreq                      : IN    STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- User DMA control for each DMA channel
  comp_done                      : IN    STD_LOGIC;
  
 --version of RBF
  rbf_version                    : IN    STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- RBF_Info[7..0]
  almost_full_wr                 : IN    STD_LOGIC;                          -- status_wr[1]
  empty_wr                       : IN    STD_LOGIC;                          -- status_wr[2]
  almost_empty_rd                : IN    STD_LOGIC;                          -- status_rd[0]
  almost_full_rd                 : IN    STD_LOGIC;                          -- status_rd[1]
  empty_rd                       : IN    STD_LOGIC;                          -- status_rd[2]
  addr_1v                        : OUT   arr_19x0_31x0;
  addr_2v                        : OUT   arr_19x0_31x0;
  addr_3v                        : OUT   arr_19x0_31x0;
  gc_and_en                      : OUT   STD_LOGIC_VECTOR( 19 DOWNTO 0 );
  R                              : OUT   arr_2x0_31x0;
  and_gt_id                      : OUT   arr_39x0_31x0;
  layer_num                      : OUT   STD_LOGIC_VECTOR( 31 DOWNTO 0 );
  addr_1v_xor                    : OUT   arr_19x0_31x0;
  addr_2v_xor                    : OUT   arr_19x0_31x0;
  addr_3v_xor                    : OUT   arr_19x0_31x0;
  gc_xor_en                      : OUT   STD_LOGIC_VECTOR( 19 DOWNTO 0 );
  xor_gt_id                      : OUT   arr_19x0_31x0;
  sel_mp_wr                      : OUT   STD_LOGIC;                          -- select for mp_wr
  sel_start_mp_wr                : OUT   STD_LOGIC;                          -- select for start_mp_wr
  sel_mp_rd                      : OUT   STD_LOGIC;                          -- select for mp_rd
  sel_start_mp_rd                : OUT   STD_LOGIC;                          -- select for start_mp_rd
  g_dreq_rd                      : IN    STD_LOGIC;                          -- Gidel DREQ signals
  g_dreq_wr                      : IN    STD_LOGIC                           -- Gidel DREQ signals
     );
 END   COMPONENT;
  
  
  
 --g_mp_pll_sv
 COMPONENT   g_mp_pll_sv
     PORT(
  clrn                           : IN    STD_LOGIC;
  mem_ref_clk                    : IN    STD_LOGIC;
  pll_mem_clk                    : OUT   STD_LOGIC;
  pll_write_clk                  : OUT   STD_LOGIC;
  pll_write_clk_pre_phy_clk      : OUT   STD_LOGIC;
  pll_addr_cmd_clk               : OUT   STD_LOGIC;
  pll_hr_clk                     : OUT   STD_LOGIC;
  pll_p2c_read_clk               : OUT   STD_LOGIC;
  pll_c2p_write_clk              : OUT   STD_LOGIC;
  pll_avl_clk                    : OUT   STD_LOGIC;
  pll_config_clk                 : OUT   STD_LOGIC;
  pll_locked                     : OUT   STD_LOGIC;
  afi_clk                        : OUT   STD_LOGIC;
  afi_half_clk                   : OUT   STD_LOGIC 
     );
 END   COMPONENT;
  
  
  
  
 COMPONENT   gc_comp
     PORT(
  
 --Internal Bus Connections
  clrn                           : IN    STD_LOGIC;                          -- 0: global reset 
  lclk                           : IN    STD_LOGIC;                          -- Clock
  addr_1v                        : IN    arr_19x0_31x0;
  addr_2v                        : IN    arr_19x0_31x0;
  addr_3v                        : IN    arr_19x0_31x0;
  comp_done                      : OUT   STD_LOGIC;
  gc_and_en                      : IN    STD_LOGIC_VECTOR( 19 DOWNTO 0 );
  R                              : IN    arr_2x0_31x0;
  and_gt_id                      : IN    arr_39x0_31x0;
  layer_num                      : IN    STD_LOGIC_VECTOR( 31 DOWNTO 0 );
  addr_1v_xor                    : IN    arr_19x0_31x0;
  addr_2v_xor                    : IN    arr_19x0_31x0;
  addr_3v_xor                    : IN    arr_19x0_31x0;
  gc_xor_en                      : IN    STD_LOGIC_VECTOR( 19 DOWNTO 0 );
  xor_gt_id                      : IN    arr_19x0_31x0;
  Bank_B_ready                   : IN    STD_LOGIC;                          -- 1: Memory controller is ready for use, 0: Initializing (due to reset)
  select_gc                      : OUT   STD_LOGIC;                          -- Port select (enable) signal. Should be high until ready comes to transfer current datatransfers data on each port clock
  data_gc_in                     : OUT   STD_LOGIC_VECTOR( 511 DOWNTO 0 );   -- Data to port gc of MultiPort mp
  data_gc_out                    : IN    STD_LOGIC_VECTOR( 511 DOWNTO 0 );   -- Data from port gc of MultiPort mp
  gc_be                          : OUT   STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Random port byte enable bits
  addr_gc                        : OUT   STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- Port address. Apply the new address to this bus before selecting the port (select=VCC)
  write_gc                       : OUT   STD_LOGIC;                          -- Port read\write signal. Assert high to write to the port
  ready_gc                       : IN    STD_LOGIC                           -- Port ready flag (goes high when the data is ready)
     );
 END   COMPONENT;
  
  
 COMPONENT   IC_1_Bank_B_Ctrl
     PORT(
  
 --Global MultiPort Connections
  clrn                           : IN    STD_LOGIC;                          -- MultiPort async global reset
  ref_clk                        : IN    STD_LOGIC;                          -- mem ref clock
  pll_mem_clk                    : IN    STD_LOGIC;
  pll_write_clk                  : IN    STD_LOGIC;
  pll_write_clk_pre_phy_clk      : IN    STD_LOGIC;
  pll_addr_cmd_clk               : IN    STD_LOGIC;
  pll_hr_clk                     : IN    STD_LOGIC;
  pll_p2c_read_clk               : IN    STD_LOGIC;
  pll_c2p_write_clk              : IN    STD_LOGIC;
  pll_avl_clk                    : IN    STD_LOGIC;
  pll_config_clk                 : IN    STD_LOGIC;
  pll_locked                     : IN    STD_LOGIC;
  afi_clk                        : IN    STD_LOGIC;
  afi_half_clk                   : IN    STD_LOGIC;
  g_reserved_control             : IN    STD_LOGIC_VECTOR( 99 DOWNTO 0 );    -- SDRAM Connection
  ready                          : OUT   STD_LOGIC;                          -- 1: Memory controller is ready for use, 0: Initializing (due to reset)
  
 --SDRAM Connections
  data                           : INOUT STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Memory data
  addr                           : OUT   STD_LOGIC_VECTOR( 15 DOWNTO 0 );    -- Memory address
  dqm                            : OUT   STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- DQM signal from MultiPort
  dqs                            : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- DQS signal from MultiPort
  dqsn                           : INOUT STD_LOGIC_VECTOR( 7  DOWNTO 0 );    -- DQSN signal from MultiPort
  ba                             : OUT   STD_LOGIC_VECTOR( 2  DOWNTO 0 );    -- SDRAM control signal
  cs_bus                         : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Chip Select signal from MultiPort
  ce                             : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- Clock Enable signal from MultiPort
  ras                            : OUT   STD_LOGIC;                          -- RAS signal from MultiPort
  cas                            : OUT   STD_LOGIC;                          -- CAS signal from MultiPort
  we                             : OUT   STD_LOGIC;                          -- Write Enable signal from MultiPort
  odt                            : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- ODT signal from MultiPort
  ck                             : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- CK
  ckn                            : OUT   STD_LOGIC_VECTOR( 1  DOWNTO 0 );    -- CKN
  oct_rzqin                      : IN    STD_LOGIC;                          -- RZK signal from MultiPort
  event_in                       : IN    STD_LOGIC;                          -- event signal from MultiPort
  mem_reset_n                    : OUT   STD_LOGIC;                          -- resetn signal from MultiPort
  
 --Port wr Connections
  clk_wr                         : IN    STD_LOGIC;                          -- Port clock
  start_wr                       : IN    STD_LOGIC;                          -- Port start (reset) signal
  select_wr                      : IN    STD_LOGIC;                          -- Port select (enable) signal
  data_wr                        : IN    STD_LOGIC_VECTOR( 255 DOWNTO 0 );   -- Data to port wr of MultiPort mp
  empty_wr                       : OUT   STD_LOGIC;                          -- Port empty flag (goes high when the internal FIFO is empty)
  almost_full_wr                 : OUT   STD_LOGIC;                          -- Port almost_full flag (goes high when the internal FIFO more than 7/8 full)
  port_error_wr                  : OUT   STD_LOGIC;                          -- Port port_error flag (goes high when an error occur to port (read from empty FIFO or write to full FIFO)
  g_dreq_mp_wr                   : OUT   STD_LOGIC;                          -- DMA transfer hold request from the port
  
 --Port rd Connections
  clk_rd                         : IN    STD_LOGIC;                          -- Port clock
  start_rd                       : IN    STD_LOGIC;                          -- Port start (reset) signal
  select_rd                      : IN    STD_LOGIC;                          -- Port select (enable) signal
  data_rd                        : OUT   STD_LOGIC_VECTOR( 255 DOWNTO 0 );   -- Data from port rd of MultiPort mp
  empty_rd                       : OUT   STD_LOGIC;                          -- Port empty flag (goes high when the internal FIFO is empty)
  almost_empty_rd                : OUT   STD_LOGIC;                          -- Port almost_empty flag (goes low when the internal FIFO more than 1/8 full)
  almost_full_rd                 : OUT   STD_LOGIC;                          -- Port almost_full flag (goes high when the internal FIFO more than 7/8 full)
  port_error_rd                  : OUT   STD_LOGIC;                          -- Port port_error flag (goes high when an error occur to port (read from empty FIFO or write to full FIFO)
  g_dreq_mp_rd                   : OUT   STD_LOGIC;                          -- DMA transfer hold request from the port
  
 --Port gc Connections
  clk_gc                         : IN    STD_LOGIC;                          -- Port clock
  select_gc                      : IN    STD_LOGIC;                          -- Port select (enable) signal
  data_gc_in                     : IN    STD_LOGIC_VECTOR( 511 DOWNTO 0 );   -- Data to port gc of MultiPort mp
  data_gc_out                    : OUT   STD_LOGIC_VECTOR( 511 DOWNTO 0 );   -- Data from port gc of MultiPort mp
  gc_be                          : IN    STD_LOGIC_VECTOR( 63 DOWNTO 0 );    -- Random port byte enable bits
  addr_gc                        : IN    STD_LOGIC_VECTOR( 31 DOWNTO 0 );    -- Port address input
  write_gc                       : IN    STD_LOGIC;                          -- Port read\write signal
  ready_gc                       : OUT   STD_LOGIC                           -- Port ready flag (goes high when the data is ready)
     );
 END   COMPONENT;
  
  
  
 --Clocks & Globals
  
 --Hardware status registers (FPGA->Host)
 SIGNAL   comp_done                  : STD_LOGIC;
 SIGNAL   rbf_version                : STD_LOGIC_VECTOR( 7  DOWNTO 0 );     -- RBF_Info[7..0]
 SIGNAL   almost_full_wr             : STD_LOGIC;                           -- status_wr[1]
 SIGNAL   empty_wr                   : STD_LOGIC;                           -- status_wr[2]
 SIGNAL   almost_empty_rd            : STD_LOGIC;                           -- status_rd[0]
 SIGNAL   almost_full_rd             : STD_LOGIC;                           -- status_rd[1]
 SIGNAL   empty_rd                   : STD_LOGIC;                           -- status_rd[2]
  
 --Mode registers (Host->FPGA). Use to set hardware working modes
 SIGNAL   clk0                       : STD_LOGIC;                           -- Main system clock, the max frequency is 300 MHZ
 SIGNAL   clk                        : STD_LOGIC;                           -- User clock, the frequency is twice/triply the frequency of clk0
 SIGNAL   clk2                       : STD_LOGIC;                           -- Is an auxiliary clock that may be used as a slow emulation clock
 SIGNAL   mem_ref_clk_int            : STD_LOGIC;                           -- Is an internal (from PLL) memory reference clock (125MHz)
 SIGNAL   id                         : STD_LOGIC_VECTOR( 2  DOWNTO 0 );     -- FPGA number identification
 SIGNAL   g_reserved_control         : STD_LOGIC_VECTOR( 99 DOWNTO 0 );     -- Gidel reserved control bus
  
 --Internal Bus Interface Signals
 SIGNAL   clrn                       : STD_LOGIC;                           -- User Global Clear   (0: clear all)
 SIGNAL   lclk                       : STD_LOGIC;                           -- Local Bus Clock
 SIGNAL   l_wr                       : STD_LOGIC;                           -- User Write Signal (1:write)
 SIGNAL   addr_wr                    : STD_LOGIC_VECTOR( 31 DOWNTO 0 );     -- local bus address for write operations
 SIGNAL   l_data_wr                  : STD_LOGIC_VECTOR( 255 DOWNTO 0 );    -- user input local data bus
 SIGNAL   mem_ready_wr               : STD_LOGIC;                           -- 1: write memory data is valid (memory is ready)
 SIGNAL   l_rd                       : STD_LOGIC;                           -- User Read Signal (0:read)
 SIGNAL   addr_rd                    : STD_LOGIC_VECTOR( 31 DOWNTO 0 );     -- local bus address for read operations
 SIGNAL   l_data_rd                  : STD_LOGIC_VECTOR( 255 DOWNTO 0 );    -- data to read back from device memories
 SIGNAL   mem_ready_rd               : STD_LOGIC;                           -- 1: end of data read transfer (memory data is valid)
  
 --User interrupt signals
 SIGNAL   interrupt                  : STD_LOGIC;                           -- Interrupt signal - assert low to send interrupt to SoftWare, when interrupt_ack is high.
 SIGNAL   interrupt_ack              : STD_LOGIC;                           -- Interrupt acknowledge signal - asserted high to to enable user interrupt.
  
 --User DREQ signals
 SIGNAL   user_dreq                  : STD_LOGIC_VECTOR( 31 DOWNTO 0 );     -- DMA control - assert low to enable DMA operation, high to stop DMA (for each DMA channel).
  
 --Other signals
 SIGNAL   addr_1v                    : arr_19x0_31x0;
 SIGNAL   addr_2v                    : arr_19x0_31x0;
 SIGNAL   addr_3v                    : arr_19x0_31x0;
 SIGNAL   gc_and_en                  : STD_LOGIC_VECTOR( 19 DOWNTO 0 );
 SIGNAL   R                          : arr_2x0_31x0;
 SIGNAL   and_gt_id                  : arr_39x0_31x0;
 SIGNAL   layer_num                  : STD_LOGIC_VECTOR( 31 DOWNTO 0 );
 SIGNAL   addr_1v_xor                : arr_19x0_31x0;
 SIGNAL   addr_2v_xor                : arr_19x0_31x0;
 SIGNAL   addr_3v_xor                : arr_19x0_31x0;
 SIGNAL   gc_xor_en                  : STD_LOGIC_VECTOR( 19 DOWNTO 0 );
 SIGNAL   xor_gt_id                  : arr_19x0_31x0;
  
 --Select signals for user's memories / reggroups
 SIGNAL   sel_mp_wr                  : STD_LOGIC;                           -- select for mp_wr
 SIGNAL   sel_start_mp_wr            : STD_LOGIC;                           -- select for start_mp_wr
 SIGNAL   sel_mp_rd                  : STD_LOGIC;                           -- select for mp_rd
 SIGNAL   sel_start_mp_rd            : STD_LOGIC;                           -- select for start_mp_rd
  
 --PROCMultiPort mp
 SIGNAL   pll_mem_clk                : STD_LOGIC;
 SIGNAL   pll_write_clk              : STD_LOGIC;
 SIGNAL   pll_write_clk_pre_phy_clk  : STD_LOGIC;
 SIGNAL   pll_addr_cmd_clk           : STD_LOGIC;
 SIGNAL   pll_hr_clk                 : STD_LOGIC;
 SIGNAL   pll_p2c_read_clk           : STD_LOGIC;
 SIGNAL   pll_c2p_write_clk          : STD_LOGIC;
 SIGNAL   pll_avl_clk                : STD_LOGIC;
 SIGNAL   pll_config_clk             : STD_LOGIC;
 SIGNAL   pll_locked                 : STD_LOGIC;
 SIGNAL   afi_clk                    : STD_LOGIC;
 SIGNAL   afi_half_clk               : STD_LOGIC;
 SIGNAL   Bank_B_ready               : STD_LOGIC;                           -- 1: Memory controller is ready for use, 0: Initializing (due to reset)
 SIGNAL   port_error_wr              : STD_LOGIC;                           -- Port port_error flag (goes high when an error occur to port (read from empty FIFO or write to full FIFO)
 SIGNAL   g_dreq_mp_wr               : STD_LOGIC;                           -- DMA transfer hold request from the port
 SIGNAL   data_rd                    : STD_LOGIC_VECTOR( 255 DOWNTO 0 );    -- Data from port rd of MultiPort mp
 SIGNAL   port_error_rd              : STD_LOGIC;                           -- Port port_error flag (goes high when an error occur to port (read from empty FIFO or write to full FIFO)
 SIGNAL   g_dreq_mp_rd               : STD_LOGIC;                           -- DMA transfer hold request from the port
 SIGNAL   select_gc                  : STD_LOGIC;                           -- Port select (enable) signal
 SIGNAL   data_gc_in                 : STD_LOGIC_VECTOR( 511 DOWNTO 0 );    -- Data to port gc of MultiPort mp
 SIGNAL   data_gc_out                : STD_LOGIC_VECTOR( 511 DOWNTO 0 );    -- Data from port gc of MultiPort mp
 SIGNAL   gc_be                      : STD_LOGIC_VECTOR( 63 DOWNTO 0 );     -- Random port byte enable bits
 SIGNAL   addr_gc                    : STD_LOGIC_VECTOR( 31 DOWNTO 0 );     -- Port address input
 SIGNAL   write_gc                   : STD_LOGIC;                           -- Port read\write signal
 SIGNAL   ready_gc                   : STD_LOGIC;                           -- Port ready flag (goes high when the data is ready)
  
  
 BEGIN
   
   
   
  --======================================================================
  --=    The Interface entity connections (connections to the host)      =
  --======================================================================
  if_dma : dma_if
  PORT MAP  (
   
  --Clocks & Globals
  ref_clk                      =>  ref_clk,                                  -- IN        25 MHz reference clock input pin
  clk0                         =>  clk0,                                     -- OUT       Main system clock, the max frequency is 300 MHZ
  clk                          =>  clk,                                      -- OUT       User clock, the frequency is twice/triply the frequency of clk0
  clk2                         =>  clk2,                                     -- OUT       Is an auxiliary clock that may be used as a slow emulation clock
  mem_ref_clk_int              =>  mem_ref_clk_int,                          -- OUT       Is an internal (from PLL) memory reference clock (125MHz)
  scl                          =>  scl,                                      -- INOUT     Serial clock. Used to synchronize communication to and from the I2C bus
  sda                          =>  sda,                                      -- INOUT     Serial data: Used to transfer addresses and data into and out of the I2C bus
  status_ledn( 3  DOWNTO 1 )   =>  status_ledn( 3  DOWNTO 1 ),               -- OUT       Status LEDs; 0: light on
  id( 2  DOWNTO 0 )            =>  id( 2  DOWNTO 0 ),                        -- OUT       FPGA number identification
  g_reserved( 33 DOWNTO 0 )    =>  g_reserved( 33 DOWNTO 0 ),                -- INOUT     Gidel reserved IO bus
  g_reserved_control( 99 DOWNTO 0 )  =>  g_reserved_control( 99 DOWNTO 0 ),  -- OUT       Gidel reserved control bus (out)
   
  --PCIe connection
  pcie_refclk                  =>  pcie_refclk,                              -- IN        Reference clock for the Hard IP for PCI Express
  pcie_perst                   =>  pcie_perst,                               -- IN        Active low reset from the PCIe reset pin of the device
  pcie_rx( 7  DOWNTO 0 )       =>  pcie_rx( 7  DOWNTO 0 ),                   -- IN        Receive inputs. These signals are the serial inputs of lanes 7�0
  pcie_tx( 7  DOWNTO 0 )       =>  pcie_tx( 7  DOWNTO 0 ),                   -- OUT       Transmit outputs. These signals are the serial outputs of lanes 7�0
   
  --Internal Bus Interface Signals
  clrn                         =>  clrn,                                     -- OUT       User Global Clear   (0: clear all)
  lclk                         =>  lclk,                                     -- OUT       Local Bus Clock
  l_wr                         =>  l_wr,                                     -- OUT       User Write Signal (1:write)
  addr_wr( 31 DOWNTO 0 )       =>  addr_wr( 31 DOWNTO 0 ),                   -- OUT       local bus address for write operations (including burst auto address increment)
  l_data_wr( 255 DOWNTO 0 )    =>  l_data_wr( 255 DOWNTO 0 ),                -- OUT       user input local data bus
  mem_ready_wr                 =>  mem_ready_wr,                             -- IN        1: end of data write transfer (memory data is valid) on rising edge of lclk
  l_rd                         =>  l_rd,                                     -- OUT       User Read Signal (0:read)
  addr_rd( 31 DOWNTO 0 )       =>  addr_rd( 31 DOWNTO 0 ),                   -- OUT       local bus address for read operations (including burst auto address increment)
  l_data_rd( 255 DOWNTO 0 )    =>  l_data_rd( 255 DOWNTO 0 ),                -- IN        data to read back from device memories
  mem_ready_rd                 =>  mem_ready_rd,                             -- IN        1: end of data read transfer (memory data is valid) on rising edge of lclk
   
  --Interrupt Logic
  interrupt                    =>  interrupt,                                -- IN        User interrupt
  interrupt_ack                =>  interrupt_ack,                            -- OUT       User interrupt acknowledge
   
  --DREQ Logic
  user_dreq( 31 DOWNTO 0 )     =>  user_dreq( 31 DOWNTO 0 ),                 -- IN        User DMA control for each DMA channel
   
  --Hardware status registers (FPGA->Host)
  comp_done                    =>  comp_done,                                -- IN   
  rbf_version( 7  DOWNTO 0 )   =>  rbf_version( 7  DOWNTO 0 ),               -- IN        RBF_Info[7..0]
  almost_full_wr               =>  almost_full_wr,                           -- IN        status_wr[1]
  empty_wr                     =>  empty_wr,                                 -- IN        status_wr[2]
  almost_empty_rd              =>  almost_empty_rd,                          -- IN        status_rd[0]
  almost_full_rd               =>  almost_full_rd,                           -- IN        status_rd[1]
  empty_rd                     =>  empty_rd,                                 -- IN        status_rd[2]
   
  --Mode registers (Host->FPGA). Use to set hardware working modes
  addr_1v                      =>  addr_1v,                                  -- OUT  
  addr_2v                      =>  addr_2v,                                  -- OUT  
  addr_3v                      =>  addr_3v,                                  -- OUT  
  gc_and_en( 19 DOWNTO 0 )     =>  gc_and_en( 19 DOWNTO 0 ),                 -- OUT  
  R                            =>  R,                                        -- OUT  
  and_gt_id                    =>  and_gt_id,                                -- OUT  
  layer_num( 31 DOWNTO 0 )     =>  layer_num( 31 DOWNTO 0 ),                 -- OUT  
  addr_1v_xor                  =>  addr_1v_xor,                              -- OUT  
  addr_2v_xor                  =>  addr_2v_xor,                              -- OUT  
  addr_3v_xor                  =>  addr_3v_xor,                              -- OUT  
  gc_xor_en( 19 DOWNTO 0 )     =>  gc_xor_en( 19 DOWNTO 0 ),                 -- OUT  
  xor_gt_id                    =>  xor_gt_id,                                -- OUT  
   
  --Select signals for user's memories / reggroups
  sel_mp_wr                    =>  sel_mp_wr,                                -- OUT       select for mp_wr
  sel_start_mp_wr              =>  sel_start_mp_wr,                          -- OUT       select for start_mp_wr
  sel_mp_rd                    =>  sel_mp_rd,                                -- OUT       select for mp_rd
  sel_start_mp_rd              =>  sel_start_mp_rd,                          -- OUT       select for start_mp_rd
  g_dreq_wr                    =>  g_dreq_mp_wr,                             -- IN   
  g_dreq_rd                    =>  g_dreq_mp_rd                              -- IN   
  );

   
   
   
  --g_mp_pll_sv
  g_mp_pll_sv_cmp : g_mp_pll_sv
  PORT MAP  (
  clrn                         =>  clrn,                                     -- IN   
  mem_ref_clk                  =>  mem_ref_clk,                              -- IN   
  pll_mem_clk                  =>  pll_mem_clk,                              -- OUT  
  pll_write_clk                =>  pll_write_clk,                            -- OUT  
  pll_write_clk_pre_phy_clk    =>  pll_write_clk_pre_phy_clk,                -- OUT  
  pll_addr_cmd_clk             =>  pll_addr_cmd_clk,                         -- OUT  
  pll_hr_clk                   =>  pll_hr_clk,                               -- OUT  
  pll_p2c_read_clk             =>  pll_p2c_read_clk,                         -- OUT  
  pll_c2p_write_clk            =>  pll_c2p_write_clk,                        -- OUT  
  pll_avl_clk                  =>  pll_avl_clk,                              -- OUT  
  pll_config_clk               =>  pll_config_clk,                           -- OUT  
  pll_locked                   =>  pll_locked,                               -- OUT  
  afi_clk                      =>  afi_clk,                                  -- OUT  
  afi_half_clk                 =>  afi_half_clk                              -- OUT  
  );

   
   
   
  --======================================================================
  --=                   User's entities' connections                     =
  --======================================================================
   
  gc_comp_cmp : gc_comp
  PORT MAP  (
  clrn                         =>  clrn,                                     -- IN   
  lclk                         =>  lclk,                                     -- IN   
  addr_1v                      =>  addr_1v,                                  -- IN   
  addr_2v                      =>  addr_2v,                                  -- IN   
  addr_3v                      =>  addr_3v,                                  -- IN   
  comp_done                    =>  comp_done,                                -- OUT  
  gc_and_en                    =>  gc_and_en,                                -- IN   
  R                            =>  R,                                        -- IN   
  and_gt_id                    =>  and_gt_id,                                -- IN   
  layer_num                    =>  layer_num,                                -- IN   
  addr_1v_xor                  =>  addr_1v_xor,                              -- IN   
  addr_2v_xor                  =>  addr_2v_xor,                              -- IN   
  addr_3v_xor                  =>  addr_3v_xor,                              -- IN   
  gc_xor_en                    =>  gc_xor_en,                                -- IN   
  xor_gt_id                    =>  xor_gt_id,                                -- IN   
  Bank_B_ready                 =>  Bank_B_ready,                             -- IN        1: Memory controller is ready for use, 0: Initializing (due to reset)
  select_gc                    =>  select_gc,                                -- OUT       Port select (enable) signal. Should be high until ready comes to transfer current datatransfers data on each port clock
  data_gc_in                   =>  data_gc_in,                               -- OUT       Data to port gc of MultiPort mp
  data_gc_out                  =>  data_gc_out,                              -- IN        Data from port gc of MultiPort mp
  gc_be                        =>  gc_be,                                    -- OUT       Random port byte enable bits
  addr_gc                      =>  addr_gc,                                  -- OUT       Port address. Apply the new address to this bus before selecting the port (select=VCC)
  write_gc                     =>  write_gc,                                 -- OUT       Port read\write signal. Assert high to write to the port
  ready_gc                     =>  ready_gc                                  -- IN        Port ready flag (goes high when the data is ready)
  );

   
   
   
   
  --======================================================================
  --=                   SDRAM controllers' connections                   =
  --======================================================================
   
  --======================================================================
  --=                         IC_1_Bank_B_Ctrl                           =
  --======================================================================
   
   
  IC_1_Bank_B_Ctrl_cmp : IC_1_Bank_B_Ctrl
  PORT MAP  (
   
  --Global MultiPort Connections
  clrn                         =>  clrn,                                     -- IN   
  ref_clk                      =>  mem_ref_clk,                              -- IN   
  pll_mem_clk                  =>  pll_mem_clk,                              -- IN   
  pll_write_clk                =>  pll_write_clk,                            -- IN   
  pll_write_clk_pre_phy_clk    =>  pll_write_clk_pre_phy_clk,                -- IN   
  pll_addr_cmd_clk             =>  pll_addr_cmd_clk,                         -- IN   
  pll_hr_clk                   =>  pll_hr_clk,                               -- IN   
  pll_p2c_read_clk             =>  pll_p2c_read_clk,                         -- IN   
  pll_c2p_write_clk            =>  pll_c2p_write_clk,                        -- IN   
  pll_avl_clk                  =>  pll_avl_clk,                              -- IN   
  pll_config_clk               =>  pll_config_clk,                           -- IN   
  pll_locked                   =>  pll_locked,                               -- IN   
  afi_clk                      =>  afi_clk,                                  -- IN   
  afi_half_clk                 =>  afi_half_clk,                             -- IN   
  g_reserved_control( 99 DOWNTO 0 )  =>  g_reserved_control( 99 DOWNTO 0 ),  -- IN   
  ready                        =>  Bank_B_ready,                             -- OUT  
   
  --SDRAM Connections
  data( 63 DOWNTO 0 )          =>  dq_b( 63 DOWNTO 0 ),                      -- OUT  
  addr( 15 DOWNTO 0 )          =>  addr_b( 15 DOWNTO 0 ),                    -- OUT  
  dqm( 7  DOWNTO 0 )           =>  dqm_b( 7  DOWNTO 0 ),                     -- OUT  
  dqs( 7  DOWNTO 0 )           =>  dqs_b( 7  DOWNTO 0 ),                     -- OUT  
  dqsn( 7  DOWNTO 0 )          =>  dqsn_b( 7  DOWNTO 0 ),                    -- OUT  
  ba( 2  DOWNTO 0 )            =>  ba_b( 2  DOWNTO 0 ),                      -- OUT  
  cs_bus( 1  DOWNTO 0 )        =>  cs_b( 1  DOWNTO 0 ),                      -- OUT  
  ce( 1  DOWNTO 0 )            =>  cke_b( 1  DOWNTO 0 ),                     -- OUT  
  ras                          =>  ras_b,                                    -- OUT  
  cas                          =>  cas_b,                                    -- OUT  
  we                           =>  we_b,                                     -- OUT  
  odt( 1  DOWNTO 0 )           =>  odt_b( 1  DOWNTO 0 ),                     -- OUT  
  ck( 1  DOWNTO 0 )            =>  ck_b( 1  DOWNTO 0 ),                      -- OUT  
  ckn( 1  DOWNTO 0 )           =>  ckn_b( 1  DOWNTO 0 ),                     -- OUT  
  oct_rzqin                    =>  rzq_b,                                    -- OUT  
  event_in                     =>  event_b,                                  -- OUT  
  mem_reset_n                  =>  resetn_b,                                 -- OUT  
   
  --Port wr Connections
  clk_wr                       =>  lclk,                                     -- IN   
  start_wr                     =>  sel_start_mp_wr,                          -- IN   
  select_wr                    =>  sel_mp_wr,                                -- IN   
  data_wr( 255 DOWNTO 0 )      =>  l_data_wr( 255 DOWNTO 0 ),                -- IN   
  empty_wr                     =>  empty_wr,                                 -- OUT  
  almost_full_wr               =>  almost_full_wr,                           -- OUT  
  port_error_wr                =>  port_error_wr,                            -- OUT  
  g_dreq_mp_wr                 =>  g_dreq_mp_wr,                             -- OUT  
   
  --Port rd Connections
  clk_rd                       =>  lclk,                                     -- IN   
  start_rd                     =>  sel_start_mp_rd,                          -- IN   
  select_rd                    =>  sel_mp_rd,                                -- IN   
  data_rd( 255 DOWNTO 0 )      =>  data_rd( 255 DOWNTO 0 ),                  -- OUT  
  empty_rd                     =>  empty_rd,                                 -- OUT  
  almost_empty_rd              =>  almost_empty_rd,                          -- OUT  
  almost_full_rd               =>  almost_full_rd,                           -- OUT  
  port_error_rd                =>  port_error_rd,                            -- OUT  
  g_dreq_mp_rd                 =>  g_dreq_mp_rd,                             -- OUT  
   
  --Port gc Connections
  clk_gc                       =>  lclk,                                     -- IN   
  select_gc                    =>  select_gc,                                -- IN   
  data_gc_in( 511 DOWNTO 0 )   =>  data_gc_in( 511 DOWNTO 0 ),               -- IN   
  data_gc_out( 511 DOWNTO 0 )  =>  data_gc_out( 511 DOWNTO 0 ),              -- OUT  
  gc_be( 63 DOWNTO 0 )         =>  gc_be( 63 DOWNTO 0 ),                     -- IN   
  addr_gc( 31 DOWNTO 0 )       =>  addr_gc( 31 DOWNTO 0 ),                   -- IN   
  write_gc                     =>  write_gc,                                 -- IN   
  ready_gc                     =>  ready_gc                                  -- OUT  
  );

   
   
  rbf_version(7 DOWNTO 0)    <=    RBF_VERSION_VAL;  
   
   
  --======================================================================
  --=                Default Values of Board Connections                 =
  --======================================================================
   
  --DDR Block C Connections
  addr_c                       <=  ( others => '0' );
  ba_c                         <=  ( others => '0' );
  cas_c                        <=  '1';
  cke_c                        <=  ( others => '0' );
  ck_c                         <=  ( others => 'Z' );
  ckn_c                        <=  ( others => 'Z' );
  cs_c                         <=  ( others => '1' );
  dq_c                         <=  ( others => 'Z' );
  dqm_c                        <=  ( others => '0' );
  dqs_c                        <=  ( others => 'Z' );
  dqsn_c                       <=  ( others => 'Z' );
  we_c                         <=  '0';
  ras_c                        <=  '1';
  odt_c                        <=  ( others => '0' );
  resetn_c                     <=  '0';
   
  --DDR Block D Connections
  dq_d                         <=  ( others => 'Z' );
  ldn_d                        <=  '1';
  bwsn_d                       <=  ( others => '0' );
  r_wn_d                       <=  '0';
  k_d                          <=  '0';
  addr_d                       <=  ( others => '0' );
   
  --DDR Block D Connections
  dq_e                         <=  ( others => 'Z' );
  ldn_e                        <=  '1';
  bwsn_e                       <=  ( others => '0' );
  r_wn_e                       <=  '0';
  k_e                          <=  '0';
  addr_e                       <=  ( others => '0' );
   
  --User's buses
   
  mem_ready_wr                 <=  '1';                                      -- '1'   NO WAIT STATES, put '0' when you want to add wait states
   
  mem_ready_rd                 <=  '1';                                      -- '1'   NO WAIT STATES, put '0' when you want to add wait states
  l_data_rd( 31 DOWNTO 0 )     <= data_rd( 31 DOWNTO 0 )   WHEN   sel_mp_rd  =  '1'   ELSE
                                ( others => '0' );
   
  l_data_rd( 255 DOWNTO 32 )   <= data_rd( 255 DOWNTO 32 )   WHEN   sel_mp_rd  =  '1'   ELSE
                                ( others => '0' );
   
  interrupt                    <=  '1';                                      -- Interrupt control - assert low to send interrupt to SoftWare, when interrupt_ack is high.
  user_dreq                    <=  ( others => '0' );                        -- DMA control - assert low to enable DMA operation, high to stop DMA (for each DMA channel).
  ledn                         <=  ( others => 'Z' );
   
  --1G PHY I/O's (Connections to on board PHY)
  phy_mdio                     <=  'Z';
  phy_mdc                      <=  '0';
  phy_resetn                   <=  '0';
  phy_tx_ctrl                  <=  '0';
  phy_tx_clk                   <=  '0';
  phy_txd                      <=  ( others => '0' );
   
  --SFP A
  sfp_link_ledn_a              <=  'Z';
  sfp_trafic_ledn_a            <=  'Z';
   
  --SFP B
  sfp_link_ledn_b              <=  'Z';
  sfp_trafic_ledn_b            <=  'Z';
   
  --L(J4) connector I/O's
  l                            <=  ( others => 'Z' );
  l_io                         <=  ( others => 'Z' );
  clk_out                      <=  ( others => '0' );
   
  --External(J3) connector I/O's
  j3_ext_io                    <=  ( others => 'Z' );
  j3_ext_io_dir                <=  ( others => '0' );                        -- Bit-0 sets direction for ext_io[7:0] and bit-1 for ext_io[11:8]. (ext_io_dir=0: Inputs, ext_io_dir=1: Outputs)
   
   
 END  dma_arch;
